`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 01/16/2025 11:06:57 PM
// Design Name: 
// Module Name: Three_One_Mux
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Three_One_Mux(
    input [31:0] a,
    input [31:0] b,
    input [31:0] c,
    output reg [31:0] out,
    input [1:0] sel
    );
    always_comb begin
        case(sel)
            2'b00: out <= a;
            2'b01: out <= b;
            2'b10: out <= c;
        endcase
    end
endmodule
